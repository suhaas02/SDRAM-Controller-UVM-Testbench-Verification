class src_sequencer extends uvm_sequencer #(transaction); 
    `uvm_component_utils(src_sequencer)

    function new(string name, uvm_component parent); 
        super.new(name, parent); 
    endfunction 

endclass