bind sdram_top checker_file assertions(.*); 